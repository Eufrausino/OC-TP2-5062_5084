module instructionMemory(
    input[31:0] readAdress,
    input clock,
    input reset,
    output[31:0] instruction
)

    

endmodule